module binding_module;
bind mem_tb mem_asserts U_assert (
.data (data),
.we (we),
.clk (clk),
.address (address),
.oe (oe),
.cs (cs)
);
endmodule